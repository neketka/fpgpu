`define MODULE_NAME fp_sub
`define SUBTRACTOR
`define NO_CE

`define MODULE_NAME fp_comp
`define NO_CE
`define AGB
`define ALB

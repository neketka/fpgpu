`define MODULE_NAME fp_sqrt
`define NO_CE

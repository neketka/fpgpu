`define MODULE_NAME fp_div
`define NO_CE
